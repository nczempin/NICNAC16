// Verilog test fixture created from schematic B:\NICNAC16\dunc16.sch - Wed Sep 17 00:13:28 2014

`timescale 1ns / 1ps

module dunc16_dunc16_sch_tb();

// Inputs
    reg CLK;
   reg RESET;

// Output
   wire I_STA;
   wire SETWRITE;
   wire CLRWRITE;
   wire WRITE;
   wire [15:0] AC_OUT;
   wire [15:0] MD_OUT;

// Bidirs

// Instantiate the UUT
   dunc16 UUT (
		.I_STA(I_STA), 
		.SETWRITE(SETWRITE), 
		.CLRWRITE(CLRWRITE), 
		.WRITE(WRITE), 
		.AC_OUT(AC_OUT), 
		.MD_OUT(MD_OUT), 
		.CLK(CLK), 
		.RESET(RESET)
   );

initial begin
CLK = 0;
	//start reset
	RESET = 1'b1;
	repeat(4)
		#10
		CLK = ~CLK;
	RESET = 1'b0;
	// end reset
	
	forever
		#10
		CLK = ~CLK; // generate a clock
end

initial begin
	@(negedge RESET); // wait for reset
	repeat (40)
	@(posedge CLK);


	$finish;
end
endmodule
